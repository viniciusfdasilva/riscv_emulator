module main

import vm

fn main() {
	vm.start_vm()
}

