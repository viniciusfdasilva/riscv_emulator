module main

import vm


mut stdin  := [1024]u8;
mut stdout := [1024]u8;


fn read(input [u8])
{

}

fn exit() {
	exit(0)
}

fn write(input [u8])
{

}

fn request_control()
{

}