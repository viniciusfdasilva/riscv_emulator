module main

import vm

fn main() {
	println('Hello World!')

	vm.start_vm()
}

